//Verilog HDL for "KALHALL_STD_LIB", "INVX1" "functional"
 
`timescale 1ns/10ps
`celldefine
module TIELO (Y);
	output Y;
	//input A;

	// Function
	buf (Y, 1'b0);

	// Timing
	specify
	endspecify
endmodule
`endcelldefine
