//Verilog HDL for "KALHALL_STD_LIB", "INVX1" "functional"
 
`timescale 1ns/10ps
`celldefine
module TIEHI (Y);
	output Y;


	// Function
	buf (Y, 1'b1);

	// Timing
	specify
	endspecify
endmodule
`endcelldefine
